// Create a module that implements a NOT gate.
module not_gate( input in, output out );
    assign out = ~in;
endmodule
